`define GIE         9'h01C
`define IER         9'h028
`define SOFTR       9'h040
`define CR 			9'h100
`define TX_FIFO 	9'h108
`define ADR 		9'h110
//`define TEN_ADR	9'h11C does not exist in my case
`define GPO			9'h124
`define TSUSTA      9'h128
`define TSUSTO      9'h12C
`define THDSTA      9'h130
`define TSUDAT      9'h134
`define TBUF 	    9'h138
`define THIGH 	    9'h13C
`define TLOW 	    9'h140
`define THDDAT 	    9'h144